`timescale 1ns / 1ps

/////////////////////////////////////////////
module ft600_mode245_tx_tb();

parameter RX_BUF_WIDTH = 4;
parameter TX_BUF_WIDTH = 4;

reg clk;
reg rst;

reg ft_clk;
wire [15:0] ft_data;
wire [1:0] ft_be;
reg ft_txe;
reg ft_rxf;
wire ft_oe;
wire ft_rd;
wire ft_wr;


initial begin
    clk = 1'b0;
    #2 // Phase
    forever #5 clk = ~clk; // 100MHz
end

initial begin
    ft_clk = 1'b0;
    // #2 // Phase
    forever #5 ft_clk = ~ft_clk; // 100MHz
end

initial begin
    rst = 1'b1;
    #1000
    rst = 1'b0;
end

reg tx_en;
reg [15:0] tx_in;
wire tx_full;

wire rx_en = 0;
wire [15:0] rx_out;
wire rx_empty;

wire tx_en2;
wire [15:0] tx_in2;

ft600_mode245 ft600(
    rst,
    clk,

    tx_en2,
    tx_in2,
    tx_full,

    rx_en,
    rx_out,
    rx_empty,

    ft_clk,
    ft_data,
    ft_be,
    ft_txe,
    ft_rxf,
    ft_oe,
    ft_rd,
    ft_wr
);

count_feeder count(
    rst,
    clk,

    tx_en2,
    tx_in2,
    tx_full
);

initial begin
    $dumpfile("ft600_mode245_tx_wave.vcd");
    $dumpvars(0, clk);
    $dumpvars(0, rst);
    $dumpvars(0, ft_clk);
    $dumpvars(0, ft_data);
    $dumpvars(0, ft_be);
    $dumpvars(0, ft_txe);
    $dumpvars(0, ft_rxf);
    $dumpvars(0, ft_oe);
    $dumpvars(0, ft_rd);
    $dumpvars(0, ft_wr);
    $dumpvars(0, tx_en);
    $dumpvars(0, tx_in);
    $dumpvars(0, tx_full);
    $dumpvars(0, rx_en);
    $dumpvars(0, rx_out);
    $dumpvars(0, rx_empty);
    $dumpvars(0, ft600);

    ft_txe = 1'b1;
    ft_rxf = 1'b1;

    tx_in = 16'hFEDC;
    tx_en = 0;

    #1200

    #10;
    tx_en = 1;
    tx_in = 16'hBEB0;

    #10;
    tx_in = 16'hBCB0;

    #10;
    tx_in = 16'hAAB0;

    #10;
    tx_en = 0;

    #10000;
    ft_txe = 0;

    #199
    ft_txe = 1;

    #100000;


    tx_in = 16'hFFAA;
    tx_en = 1;

    #10;
    tx_en = 0;

    #50
    ft_txe = 0;

    #50000;

    $finish;
end
endmodule
